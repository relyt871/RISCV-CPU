`include "def.v"

module cdb (
    //input from register
    //input from robuffer
    //output to robuffer
    //input from alu
    //output to reservationstation
    //output to lsbuffer
);

endmodule